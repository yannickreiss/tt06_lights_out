/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`define default_netname none

module tt_um_yannickreiss_lights_out (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // will go high when the design is enabled
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // All output pins must be assigned. If not used, assign to 0.
  assign uio_oe  = 8'b00000010;

  // Matrix (input)
  wire in1;
  wire in2;
  wire in3;
  wire in4;
  wire in5;
  wire in6;
  wire in7;
  wire in8;
  wire in9;
  assign in1 = ui_in[0];
  assign in2 = ui_in[1];
  assign in3 = ui_in[2];
  assign in4 = ui_in[3];
  assign in5 = ui_in[4];
  assign in6 = ui_in[5];
  assign in7 = ui_in[6];
  assign in8 = ui_in[7];
  assign in9 = uio_in[0];

  // Matrix (current field)
  reg field1;
  reg field2;
  reg field3;
  reg field4;
  reg field5;
  reg field6;
  reg field7;
  reg field8;
  reg field9;

  // Matrix (output)
  assign uo_out[0] = field1;
  assign uo_out[1] = field2;
  assign uo_out[2] = field3;
  assign uo_out[3] = field4;
  assign uo_out[4] = field5;
  assign uo_out[5] = field6;
  assign uo_out[6] = field7;
  assign uo_out[7] = field8;
  assign uio_out[0] = field9;

  // uio_out map to zero
  assign uio_out[7:1] = 7'b0;

  always @(posedge clk) begin
    if (ena == 1'b1) begin
      if (rst_n == 1'b1) begin

        // Do act normal

      end
      else begin

        // set new matrix in a pseudo random way
        field1 <= 1'b0;
        field2 <= 1'b0;
        field3 <= 1'b0;
        field4 <= 1'b0;
        field5 <= 1'b1;
        field6 <= 1'b0;
        field7 <= 1'b0;
        field8 <= 1'b0;
      end
    end
  end

endmodule
